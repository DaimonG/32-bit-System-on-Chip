##
## LEF for PtnCells ;
## created by Innovus v18.10-p002_1 on Tue Apr 20 18:55:30 2021
##

VERSION 5.5 ;

NAMESCASESENSITIVE ON ;
BUSBITCHARS "[]" ;
DIVIDERCHAR "/" ;

MACRO ensc450
  CLASS BLOCK ;
  SIZE 630.040000 BY 480.060000 ;
  FOREIGN ensc450 0.000000 0.000000 ;
  ORIGIN 0 0 ;
  SYMMETRY X Y R90 ;
  PIN clk
    DIRECTION INPUT ;
    USE SIGNAL ;
  END clk
  PIN resetn
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal2 ;
        RECT 282.970000 479.990000 283.040000 480.060000 ;
    END
  END resetn
  PIN EXT_NREADY
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal2 ;
        RECT 345.480000 0.000000 345.550000 0.070000 ;
    END
  END EXT_NREADY
  PIN EXT_BUSY
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal2 ;
        RECT 283.920000 479.990000 283.990000 480.060000 ;
    END
  END EXT_BUSY
  PIN EXT_MR
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal2 ;
        RECT 284.870000 479.990000 284.940000 480.060000 ;
    END
  END EXT_MR
  PIN EXT_MW
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal2 ;
        RECT 285.820000 479.990000 285.890000 480.060000 ;
    END
  END EXT_MW
  PIN EXT_ADDRBUS[31]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal2 ;
        RECT 316.220000 479.990000 316.290000 480.060000 ;
    END
  END EXT_ADDRBUS[31]
  PIN EXT_ADDRBUS[30]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal2 ;
        RECT 315.270000 479.990000 315.340000 480.060000 ;
    END
  END EXT_ADDRBUS[30]
  PIN EXT_ADDRBUS[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal2 ;
        RECT 314.320000 479.990000 314.390000 480.060000 ;
    END
  END EXT_ADDRBUS[29]
  PIN EXT_ADDRBUS[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal2 ;
        RECT 313.370000 479.990000 313.440000 480.060000 ;
    END
  END EXT_ADDRBUS[28]
  PIN EXT_ADDRBUS[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal2 ;
        RECT 312.420000 479.990000 312.490000 480.060000 ;
    END
  END EXT_ADDRBUS[27]
  PIN EXT_ADDRBUS[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal2 ;
        RECT 311.470000 479.990000 311.540000 480.060000 ;
    END
  END EXT_ADDRBUS[26]
  PIN EXT_ADDRBUS[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal2 ;
        RECT 310.520000 479.990000 310.590000 480.060000 ;
    END
  END EXT_ADDRBUS[25]
  PIN EXT_ADDRBUS[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal2 ;
        RECT 309.570000 479.990000 309.640000 480.060000 ;
    END
  END EXT_ADDRBUS[24]
  PIN EXT_ADDRBUS[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal2 ;
        RECT 308.620000 479.990000 308.690000 480.060000 ;
    END
  END EXT_ADDRBUS[23]
  PIN EXT_ADDRBUS[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal2 ;
        RECT 307.670000 479.990000 307.740000 480.060000 ;
    END
  END EXT_ADDRBUS[22]
  PIN EXT_ADDRBUS[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal2 ;
        RECT 306.720000 479.990000 306.790000 480.060000 ;
    END
  END EXT_ADDRBUS[21]
  PIN EXT_ADDRBUS[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal2 ;
        RECT 305.770000 479.990000 305.840000 480.060000 ;
    END
  END EXT_ADDRBUS[20]
  PIN EXT_ADDRBUS[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal2 ;
        RECT 304.820000 479.990000 304.890000 480.060000 ;
    END
  END EXT_ADDRBUS[19]
  PIN EXT_ADDRBUS[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal2 ;
        RECT 303.870000 479.990000 303.940000 480.060000 ;
    END
  END EXT_ADDRBUS[18]
  PIN EXT_ADDRBUS[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal2 ;
        RECT 302.920000 479.990000 302.990000 480.060000 ;
    END
  END EXT_ADDRBUS[17]
  PIN EXT_ADDRBUS[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal2 ;
        RECT 301.970000 479.990000 302.040000 480.060000 ;
    END
  END EXT_ADDRBUS[16]
  PIN EXT_ADDRBUS[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal2 ;
        RECT 301.020000 479.990000 301.090000 480.060000 ;
    END
  END EXT_ADDRBUS[15]
  PIN EXT_ADDRBUS[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal2 ;
        RECT 300.070000 479.990000 300.140000 480.060000 ;
    END
  END EXT_ADDRBUS[14]
  PIN EXT_ADDRBUS[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal2 ;
        RECT 299.120000 479.990000 299.190000 480.060000 ;
    END
  END EXT_ADDRBUS[13]
  PIN EXT_ADDRBUS[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal2 ;
        RECT 298.170000 479.990000 298.240000 480.060000 ;
    END
  END EXT_ADDRBUS[12]
  PIN EXT_ADDRBUS[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal2 ;
        RECT 297.220000 479.990000 297.290000 480.060000 ;
    END
  END EXT_ADDRBUS[11]
  PIN EXT_ADDRBUS[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal2 ;
        RECT 296.270000 479.990000 296.340000 480.060000 ;
    END
  END EXT_ADDRBUS[10]
  PIN EXT_ADDRBUS[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal2 ;
        RECT 295.320000 479.990000 295.390000 480.060000 ;
    END
  END EXT_ADDRBUS[9]
  PIN EXT_ADDRBUS[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal2 ;
        RECT 294.370000 479.990000 294.440000 480.060000 ;
    END
  END EXT_ADDRBUS[8]
  PIN EXT_ADDRBUS[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal2 ;
        RECT 293.420000 479.990000 293.490000 480.060000 ;
    END
  END EXT_ADDRBUS[7]
  PIN EXT_ADDRBUS[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal2 ;
        RECT 292.470000 479.990000 292.540000 480.060000 ;
    END
  END EXT_ADDRBUS[6]
  PIN EXT_ADDRBUS[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal2 ;
        RECT 291.520000 479.990000 291.590000 480.060000 ;
    END
  END EXT_ADDRBUS[5]
  PIN EXT_ADDRBUS[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal2 ;
        RECT 290.570000 479.990000 290.640000 480.060000 ;
    END
  END EXT_ADDRBUS[4]
  PIN EXT_ADDRBUS[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal2 ;
        RECT 289.620000 479.990000 289.690000 480.060000 ;
    END
  END EXT_ADDRBUS[3]
  PIN EXT_ADDRBUS[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal2 ;
        RECT 288.670000 479.990000 288.740000 480.060000 ;
    END
  END EXT_ADDRBUS[2]
  PIN EXT_ADDRBUS[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal2 ;
        RECT 287.720000 479.990000 287.790000 480.060000 ;
    END
  END EXT_ADDRBUS[1]
  PIN EXT_ADDRBUS[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal2 ;
        RECT 286.770000 479.990000 286.840000 480.060000 ;
    END
  END EXT_ADDRBUS[0]
  PIN EXT_RDATABUS[31]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal2 ;
        RECT 284.680000 0.000000 284.750000 0.070000 ;
    END
  END EXT_RDATABUS[31]
  PIN EXT_RDATABUS[30]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal2 ;
        RECT 286.580000 0.000000 286.650000 0.070000 ;
    END
  END EXT_RDATABUS[30]
  PIN EXT_RDATABUS[29]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal2 ;
        RECT 288.480000 0.000000 288.550000 0.070000 ;
    END
  END EXT_RDATABUS[29]
  PIN EXT_RDATABUS[28]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal2 ;
        RECT 290.380000 0.000000 290.450000 0.070000 ;
    END
  END EXT_RDATABUS[28]
  PIN EXT_RDATABUS[27]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal2 ;
        RECT 292.280000 0.000000 292.350000 0.070000 ;
    END
  END EXT_RDATABUS[27]
  PIN EXT_RDATABUS[26]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal2 ;
        RECT 294.180000 0.000000 294.250000 0.070000 ;
    END
  END EXT_RDATABUS[26]
  PIN EXT_RDATABUS[25]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal2 ;
        RECT 296.080000 0.000000 296.150000 0.070000 ;
    END
  END EXT_RDATABUS[25]
  PIN EXT_RDATABUS[24]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal2 ;
        RECT 297.980000 0.000000 298.050000 0.070000 ;
    END
  END EXT_RDATABUS[24]
  PIN EXT_RDATABUS[23]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal2 ;
        RECT 299.880000 0.000000 299.950000 0.070000 ;
    END
  END EXT_RDATABUS[23]
  PIN EXT_RDATABUS[22]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal2 ;
        RECT 301.780000 0.000000 301.850000 0.070000 ;
    END
  END EXT_RDATABUS[22]
  PIN EXT_RDATABUS[21]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal2 ;
        RECT 303.680000 0.000000 303.750000 0.070000 ;
    END
  END EXT_RDATABUS[21]
  PIN EXT_RDATABUS[20]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal2 ;
        RECT 305.580000 0.000000 305.650000 0.070000 ;
    END
  END EXT_RDATABUS[20]
  PIN EXT_RDATABUS[19]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal2 ;
        RECT 307.480000 0.000000 307.550000 0.070000 ;
    END
  END EXT_RDATABUS[19]
  PIN EXT_RDATABUS[18]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal2 ;
        RECT 309.380000 0.000000 309.450000 0.070000 ;
    END
  END EXT_RDATABUS[18]
  PIN EXT_RDATABUS[17]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal2 ;
        RECT 311.280000 0.000000 311.350000 0.070000 ;
    END
  END EXT_RDATABUS[17]
  PIN EXT_RDATABUS[16]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal2 ;
        RECT 313.180000 0.000000 313.250000 0.070000 ;
    END
  END EXT_RDATABUS[16]
  PIN EXT_RDATABUS[15]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal2 ;
        RECT 315.080000 0.000000 315.150000 0.070000 ;
    END
  END EXT_RDATABUS[15]
  PIN EXT_RDATABUS[14]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal2 ;
        RECT 316.980000 0.000000 317.050000 0.070000 ;
    END
  END EXT_RDATABUS[14]
  PIN EXT_RDATABUS[13]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal2 ;
        RECT 318.880000 0.000000 318.950000 0.070000 ;
    END
  END EXT_RDATABUS[13]
  PIN EXT_RDATABUS[12]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal2 ;
        RECT 320.780000 0.000000 320.850000 0.070000 ;
    END
  END EXT_RDATABUS[12]
  PIN EXT_RDATABUS[11]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal2 ;
        RECT 322.680000 0.000000 322.750000 0.070000 ;
    END
  END EXT_RDATABUS[11]
  PIN EXT_RDATABUS[10]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal2 ;
        RECT 324.580000 0.000000 324.650000 0.070000 ;
    END
  END EXT_RDATABUS[10]
  PIN EXT_RDATABUS[9]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal2 ;
        RECT 326.480000 0.000000 326.550000 0.070000 ;
    END
  END EXT_RDATABUS[9]
  PIN EXT_RDATABUS[8]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal2 ;
        RECT 328.380000 0.000000 328.450000 0.070000 ;
    END
  END EXT_RDATABUS[8]
  PIN EXT_RDATABUS[7]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal2 ;
        RECT 330.280000 0.000000 330.350000 0.070000 ;
    END
  END EXT_RDATABUS[7]
  PIN EXT_RDATABUS[6]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal2 ;
        RECT 332.180000 0.000000 332.250000 0.070000 ;
    END
  END EXT_RDATABUS[6]
  PIN EXT_RDATABUS[5]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal2 ;
        RECT 334.080000 0.000000 334.150000 0.070000 ;
    END
  END EXT_RDATABUS[5]
  PIN EXT_RDATABUS[4]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal2 ;
        RECT 335.980000 0.000000 336.050000 0.070000 ;
    END
  END EXT_RDATABUS[4]
  PIN EXT_RDATABUS[3]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal2 ;
        RECT 337.880000 0.000000 337.950000 0.070000 ;
    END
  END EXT_RDATABUS[3]
  PIN EXT_RDATABUS[2]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal2 ;
        RECT 339.780000 0.000000 339.850000 0.070000 ;
    END
  END EXT_RDATABUS[2]
  PIN EXT_RDATABUS[1]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal2 ;
        RECT 341.680000 0.000000 341.750000 0.070000 ;
    END
  END EXT_RDATABUS[1]
  PIN EXT_RDATABUS[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal2 ;
        RECT 343.580000 0.000000 343.650000 0.070000 ;
    END
  END EXT_RDATABUS[0]
  PIN EXT_WDATABUS[31]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal2 ;
        RECT 346.620000 479.990000 346.690000 480.060000 ;
    END
  END EXT_WDATABUS[31]
  PIN EXT_WDATABUS[30]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal2 ;
        RECT 345.670000 479.990000 345.740000 480.060000 ;
    END
  END EXT_WDATABUS[30]
  PIN EXT_WDATABUS[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal2 ;
        RECT 344.720000 479.990000 344.790000 480.060000 ;
    END
  END EXT_WDATABUS[29]
  PIN EXT_WDATABUS[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal2 ;
        RECT 343.770000 479.990000 343.840000 480.060000 ;
    END
  END EXT_WDATABUS[28]
  PIN EXT_WDATABUS[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal2 ;
        RECT 342.820000 479.990000 342.890000 480.060000 ;
    END
  END EXT_WDATABUS[27]
  PIN EXT_WDATABUS[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal2 ;
        RECT 341.870000 479.990000 341.940000 480.060000 ;
    END
  END EXT_WDATABUS[26]
  PIN EXT_WDATABUS[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal2 ;
        RECT 340.920000 479.990000 340.990000 480.060000 ;
    END
  END EXT_WDATABUS[25]
  PIN EXT_WDATABUS[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal2 ;
        RECT 339.970000 479.990000 340.040000 480.060000 ;
    END
  END EXT_WDATABUS[24]
  PIN EXT_WDATABUS[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal2 ;
        RECT 339.020000 479.990000 339.090000 480.060000 ;
    END
  END EXT_WDATABUS[23]
  PIN EXT_WDATABUS[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal2 ;
        RECT 338.070000 479.990000 338.140000 480.060000 ;
    END
  END EXT_WDATABUS[22]
  PIN EXT_WDATABUS[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal2 ;
        RECT 337.120000 479.990000 337.190000 480.060000 ;
    END
  END EXT_WDATABUS[21]
  PIN EXT_WDATABUS[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal2 ;
        RECT 336.170000 479.990000 336.240000 480.060000 ;
    END
  END EXT_WDATABUS[20]
  PIN EXT_WDATABUS[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal2 ;
        RECT 335.220000 479.990000 335.290000 480.060000 ;
    END
  END EXT_WDATABUS[19]
  PIN EXT_WDATABUS[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal2 ;
        RECT 334.270000 479.990000 334.340000 480.060000 ;
    END
  END EXT_WDATABUS[18]
  PIN EXT_WDATABUS[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal2 ;
        RECT 333.320000 479.990000 333.390000 480.060000 ;
    END
  END EXT_WDATABUS[17]
  PIN EXT_WDATABUS[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal2 ;
        RECT 332.370000 479.990000 332.440000 480.060000 ;
    END
  END EXT_WDATABUS[16]
  PIN EXT_WDATABUS[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal2 ;
        RECT 331.420000 479.990000 331.490000 480.060000 ;
    END
  END EXT_WDATABUS[15]
  PIN EXT_WDATABUS[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal2 ;
        RECT 330.470000 479.990000 330.540000 480.060000 ;
    END
  END EXT_WDATABUS[14]
  PIN EXT_WDATABUS[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal2 ;
        RECT 329.520000 479.990000 329.590000 480.060000 ;
    END
  END EXT_WDATABUS[13]
  PIN EXT_WDATABUS[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal2 ;
        RECT 328.570000 479.990000 328.640000 480.060000 ;
    END
  END EXT_WDATABUS[12]
  PIN EXT_WDATABUS[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal2 ;
        RECT 327.620000 479.990000 327.690000 480.060000 ;
    END
  END EXT_WDATABUS[11]
  PIN EXT_WDATABUS[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal2 ;
        RECT 326.670000 479.990000 326.740000 480.060000 ;
    END
  END EXT_WDATABUS[10]
  PIN EXT_WDATABUS[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal2 ;
        RECT 325.720000 479.990000 325.790000 480.060000 ;
    END
  END EXT_WDATABUS[9]
  PIN EXT_WDATABUS[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal2 ;
        RECT 324.770000 479.990000 324.840000 480.060000 ;
    END
  END EXT_WDATABUS[8]
  PIN EXT_WDATABUS[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal2 ;
        RECT 323.820000 479.990000 323.890000 480.060000 ;
    END
  END EXT_WDATABUS[7]
  PIN EXT_WDATABUS[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal2 ;
        RECT 322.870000 479.990000 322.940000 480.060000 ;
    END
  END EXT_WDATABUS[6]
  PIN EXT_WDATABUS[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal2 ;
        RECT 321.920000 479.990000 321.990000 480.060000 ;
    END
  END EXT_WDATABUS[5]
  PIN EXT_WDATABUS[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal2 ;
        RECT 320.970000 479.990000 321.040000 480.060000 ;
    END
  END EXT_WDATABUS[4]
  PIN EXT_WDATABUS[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal2 ;
        RECT 320.020000 479.990000 320.090000 480.060000 ;
    END
  END EXT_WDATABUS[3]
  PIN EXT_WDATABUS[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal2 ;
        RECT 319.070000 479.990000 319.140000 480.060000 ;
    END
  END EXT_WDATABUS[2]
  PIN EXT_WDATABUS[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal2 ;
        RECT 318.120000 479.990000 318.190000 480.060000 ;
    END
  END EXT_WDATABUS[1]
  PIN EXT_WDATABUS[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal2 ;
        RECT 317.170000 479.990000 317.240000 480.060000 ;
    END
  END EXT_WDATABUS[0]
  OBS
    LAYER metal1 ;
      RECT 0.000000 0.000000 630.040000 480.060000 ;
    LAYER metal2 ;
      RECT 346.760000 479.920000 630.040000 480.060000 ;
      RECT 345.810000 479.920000 346.550000 480.060000 ;
      RECT 344.860000 479.920000 345.600000 480.060000 ;
      RECT 343.910000 479.920000 344.650000 480.060000 ;
      RECT 342.960000 479.920000 343.700000 480.060000 ;
      RECT 342.010000 479.920000 342.750000 480.060000 ;
      RECT 341.060000 479.920000 341.800000 480.060000 ;
      RECT 340.110000 479.920000 340.850000 480.060000 ;
      RECT 339.160000 479.920000 339.900000 480.060000 ;
      RECT 338.210000 479.920000 338.950000 480.060000 ;
      RECT 337.260000 479.920000 338.000000 480.060000 ;
      RECT 336.310000 479.920000 337.050000 480.060000 ;
      RECT 335.360000 479.920000 336.100000 480.060000 ;
      RECT 334.410000 479.920000 335.150000 480.060000 ;
      RECT 333.460000 479.920000 334.200000 480.060000 ;
      RECT 332.510000 479.920000 333.250000 480.060000 ;
      RECT 331.560000 479.920000 332.300000 480.060000 ;
      RECT 330.610000 479.920000 331.350000 480.060000 ;
      RECT 329.660000 479.920000 330.400000 480.060000 ;
      RECT 328.710000 479.920000 329.450000 480.060000 ;
      RECT 327.760000 479.920000 328.500000 480.060000 ;
      RECT 326.810000 479.920000 327.550000 480.060000 ;
      RECT 325.860000 479.920000 326.600000 480.060000 ;
      RECT 324.910000 479.920000 325.650000 480.060000 ;
      RECT 323.960000 479.920000 324.700000 480.060000 ;
      RECT 323.010000 479.920000 323.750000 480.060000 ;
      RECT 322.060000 479.920000 322.800000 480.060000 ;
      RECT 321.110000 479.920000 321.850000 480.060000 ;
      RECT 320.160000 479.920000 320.900000 480.060000 ;
      RECT 319.210000 479.920000 319.950000 480.060000 ;
      RECT 318.260000 479.920000 319.000000 480.060000 ;
      RECT 317.310000 479.920000 318.050000 480.060000 ;
      RECT 316.360000 479.920000 317.100000 480.060000 ;
      RECT 315.410000 479.920000 316.150000 480.060000 ;
      RECT 314.460000 479.920000 315.200000 480.060000 ;
      RECT 313.510000 479.920000 314.250000 480.060000 ;
      RECT 312.560000 479.920000 313.300000 480.060000 ;
      RECT 311.610000 479.920000 312.350000 480.060000 ;
      RECT 310.660000 479.920000 311.400000 480.060000 ;
      RECT 309.710000 479.920000 310.450000 480.060000 ;
      RECT 308.760000 479.920000 309.500000 480.060000 ;
      RECT 307.810000 479.920000 308.550000 480.060000 ;
      RECT 306.860000 479.920000 307.600000 480.060000 ;
      RECT 305.910000 479.920000 306.650000 480.060000 ;
      RECT 304.960000 479.920000 305.700000 480.060000 ;
      RECT 304.010000 479.920000 304.750000 480.060000 ;
      RECT 303.060000 479.920000 303.800000 480.060000 ;
      RECT 302.110000 479.920000 302.850000 480.060000 ;
      RECT 301.160000 479.920000 301.900000 480.060000 ;
      RECT 300.210000 479.920000 300.950000 480.060000 ;
      RECT 299.260000 479.920000 300.000000 480.060000 ;
      RECT 298.310000 479.920000 299.050000 480.060000 ;
      RECT 297.360000 479.920000 298.100000 480.060000 ;
      RECT 296.410000 479.920000 297.150000 480.060000 ;
      RECT 295.460000 479.920000 296.200000 480.060000 ;
      RECT 294.510000 479.920000 295.250000 480.060000 ;
      RECT 293.560000 479.920000 294.300000 480.060000 ;
      RECT 292.610000 479.920000 293.350000 480.060000 ;
      RECT 291.660000 479.920000 292.400000 480.060000 ;
      RECT 290.710000 479.920000 291.450000 480.060000 ;
      RECT 289.760000 479.920000 290.500000 480.060000 ;
      RECT 288.810000 479.920000 289.550000 480.060000 ;
      RECT 287.860000 479.920000 288.600000 480.060000 ;
      RECT 286.910000 479.920000 287.650000 480.060000 ;
      RECT 285.960000 479.920000 286.700000 480.060000 ;
      RECT 285.010000 479.920000 285.750000 480.060000 ;
      RECT 284.060000 479.920000 284.800000 480.060000 ;
      RECT 283.110000 479.920000 283.850000 480.060000 ;
      RECT 0.000000 479.920000 282.900000 480.060000 ;
      RECT 0.000000 0.140000 630.040000 479.920000 ;
      RECT 345.620000 0.000000 630.040000 0.140000 ;
      RECT 343.720000 0.000000 345.410000 0.140000 ;
      RECT 341.820000 0.000000 343.510000 0.140000 ;
      RECT 339.920000 0.000000 341.610000 0.140000 ;
      RECT 338.020000 0.000000 339.710000 0.140000 ;
      RECT 336.120000 0.000000 337.810000 0.140000 ;
      RECT 334.220000 0.000000 335.910000 0.140000 ;
      RECT 332.320000 0.000000 334.010000 0.140000 ;
      RECT 330.420000 0.000000 332.110000 0.140000 ;
      RECT 328.520000 0.000000 330.210000 0.140000 ;
      RECT 326.620000 0.000000 328.310000 0.140000 ;
      RECT 324.720000 0.000000 326.410000 0.140000 ;
      RECT 322.820000 0.000000 324.510000 0.140000 ;
      RECT 320.920000 0.000000 322.610000 0.140000 ;
      RECT 319.020000 0.000000 320.710000 0.140000 ;
      RECT 317.120000 0.000000 318.810000 0.140000 ;
      RECT 315.220000 0.000000 316.910000 0.140000 ;
      RECT 313.320000 0.000000 315.010000 0.140000 ;
      RECT 311.420000 0.000000 313.110000 0.140000 ;
      RECT 309.520000 0.000000 311.210000 0.140000 ;
      RECT 307.620000 0.000000 309.310000 0.140000 ;
      RECT 305.720000 0.000000 307.410000 0.140000 ;
      RECT 303.820000 0.000000 305.510000 0.140000 ;
      RECT 301.920000 0.000000 303.610000 0.140000 ;
      RECT 300.020000 0.000000 301.710000 0.140000 ;
      RECT 298.120000 0.000000 299.810000 0.140000 ;
      RECT 296.220000 0.000000 297.910000 0.140000 ;
      RECT 294.320000 0.000000 296.010000 0.140000 ;
      RECT 292.420000 0.000000 294.110000 0.140000 ;
      RECT 290.520000 0.000000 292.210000 0.140000 ;
      RECT 288.620000 0.000000 290.310000 0.140000 ;
      RECT 286.720000 0.000000 288.410000 0.140000 ;
      RECT 284.820000 0.000000 286.510000 0.140000 ;
      RECT 0.000000 0.000000 284.610000 0.140000 ;
    LAYER metal3 ;
      RECT 0.000000 0.000000 630.040000 480.060000 ;
    LAYER metal4 ;
      RECT 0.000000 0.000000 630.040000 480.060000 ;
    LAYER metal5 ;
      RECT 0.000000 0.000000 630.040000 480.060000 ;
    LAYER metal6 ;
      RECT 0.000000 0.000000 630.040000 480.060000 ;
    LAYER metal7 ;
      RECT 0.000000 0.000000 630.040000 480.060000 ;
    LAYER metal8 ;
      RECT 0.000000 0.000000 630.040000 480.060000 ;
    LAYER metal9 ;
      RECT 0.000000 0.000000 630.040000 480.060000 ;
    LAYER metal10 ;
      RECT 0.000000 0.000000 630.040000 480.060000 ;
  END
END ensc450

END LIBRARY
