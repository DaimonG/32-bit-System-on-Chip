##
## LEF for PtnCells ;
## created by Innovus v18.10-p002_1 on Tue Apr 20 17:40:23 2021
##

VERSION 5.5 ;

NAMESCASESENSITIVE ON ;
BUSBITCHARS "[]" ;
DIVIDERCHAR "/" ;

MACRO aes128keyWrapper
  CLASS BLOCK ;
  SIZE 184.680000 BY 183.120000 ;
  FOREIGN aes128keyWrapper 0.000000 0.000000 ;
  ORIGIN 0 0 ;
  SYMMETRY X Y R90 ;
  PIN reset
    DIRECTION INPUT ;
    USE SIGNAL ;
  END reset
  PIN clock
    DIRECTION INPUT ;
    USE SIGNAL ;
  END clock
  PIN input[31]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal2 ;
        RECT 90.690000 183.050000 90.760000 183.120000 ;
    END
  END input[31]
  PIN input[30]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal2 ;
        RECT 89.740000 183.050000 89.810000 183.120000 ;
    END
  END input[30]
  PIN input[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal2 ;
        RECT 88.790000 183.050000 88.860000 183.120000 ;
    END
  END input[29]
  PIN input[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal2 ;
        RECT 87.840000 183.050000 87.910000 183.120000 ;
    END
  END input[28]
  PIN input[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal2 ;
        RECT 86.890000 183.050000 86.960000 183.120000 ;
    END
  END input[27]
  PIN input[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal2 ;
        RECT 85.940000 183.050000 86.010000 183.120000 ;
    END
  END input[26]
  PIN input[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal2 ;
        RECT 84.990000 183.050000 85.060000 183.120000 ;
    END
  END input[25]
  PIN input[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal2 ;
        RECT 84.040000 183.050000 84.110000 183.120000 ;
    END
  END input[24]
  PIN input[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal2 ;
        RECT 83.090000 183.050000 83.160000 183.120000 ;
    END
  END input[23]
  PIN input[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal2 ;
        RECT 82.140000 183.050000 82.210000 183.120000 ;
    END
  END input[22]
  PIN input[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal2 ;
        RECT 81.190000 183.050000 81.260000 183.120000 ;
    END
  END input[21]
  PIN input[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal2 ;
        RECT 80.240000 183.050000 80.310000 183.120000 ;
    END
  END input[20]
  PIN input[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal2 ;
        RECT 79.290000 183.050000 79.360000 183.120000 ;
    END
  END input[19]
  PIN input[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal2 ;
        RECT 78.340000 183.050000 78.410000 183.120000 ;
    END
  END input[18]
  PIN input[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal2 ;
        RECT 77.390000 183.050000 77.460000 183.120000 ;
    END
  END input[17]
  PIN input[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal2 ;
        RECT 76.440000 183.050000 76.510000 183.120000 ;
    END
  END input[16]
  PIN input[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal2 ;
        RECT 75.490000 183.050000 75.560000 183.120000 ;
    END
  END input[15]
  PIN input[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal2 ;
        RECT 74.540000 183.050000 74.610000 183.120000 ;
    END
  END input[14]
  PIN input[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal2 ;
        RECT 73.590000 183.050000 73.660000 183.120000 ;
    END
  END input[13]
  PIN input[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal2 ;
        RECT 72.640000 183.050000 72.710000 183.120000 ;
    END
  END input[12]
  PIN input[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal2 ;
        RECT 71.690000 183.050000 71.760000 183.120000 ;
    END
  END input[11]
  PIN input[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal2 ;
        RECT 70.740000 183.050000 70.810000 183.120000 ;
    END
  END input[10]
  PIN input[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal2 ;
        RECT 69.790000 183.050000 69.860000 183.120000 ;
    END
  END input[9]
  PIN input[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal2 ;
        RECT 68.840000 183.050000 68.910000 183.120000 ;
    END
  END input[8]
  PIN input[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal2 ;
        RECT 67.890000 183.050000 67.960000 183.120000 ;
    END
  END input[7]
  PIN input[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal2 ;
        RECT 66.940000 183.050000 67.010000 183.120000 ;
    END
  END input[6]
  PIN input[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal2 ;
        RECT 65.990000 183.050000 66.060000 183.120000 ;
    END
  END input[5]
  PIN input[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal2 ;
        RECT 65.040000 183.050000 65.110000 183.120000 ;
    END
  END input[4]
  PIN input[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal2 ;
        RECT 64.090000 183.050000 64.160000 183.120000 ;
    END
  END input[3]
  PIN input[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal2 ;
        RECT 63.140000 183.050000 63.210000 183.120000 ;
    END
  END input[2]
  PIN input[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal2 ;
        RECT 62.190000 183.050000 62.260000 183.120000 ;
    END
  END input[1]
  PIN input[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal2 ;
        RECT 61.240000 183.050000 61.310000 183.120000 ;
    END
  END input[0]
  PIN cipher[31]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal2 ;
        RECT 62.950000 0.000000 63.020000 0.070000 ;
    END
  END cipher[31]
  PIN cipher[30]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal2 ;
        RECT 64.850000 0.000000 64.920000 0.070000 ;
    END
  END cipher[30]
  PIN cipher[29]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal2 ;
        RECT 66.750000 0.000000 66.820000 0.070000 ;
    END
  END cipher[29]
  PIN cipher[28]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal2 ;
        RECT 68.650000 0.000000 68.720000 0.070000 ;
    END
  END cipher[28]
  PIN cipher[27]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal2 ;
        RECT 70.550000 0.000000 70.620000 0.070000 ;
    END
  END cipher[27]
  PIN cipher[26]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal2 ;
        RECT 72.450000 0.000000 72.520000 0.070000 ;
    END
  END cipher[26]
  PIN cipher[25]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal2 ;
        RECT 74.350000 0.000000 74.420000 0.070000 ;
    END
  END cipher[25]
  PIN cipher[24]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal2 ;
        RECT 76.250000 0.000000 76.320000 0.070000 ;
    END
  END cipher[24]
  PIN cipher[23]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal2 ;
        RECT 78.150000 0.000000 78.220000 0.070000 ;
    END
  END cipher[23]
  PIN cipher[22]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal2 ;
        RECT 80.050000 0.000000 80.120000 0.070000 ;
    END
  END cipher[22]
  PIN cipher[21]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal2 ;
        RECT 81.950000 0.000000 82.020000 0.070000 ;
    END
  END cipher[21]
  PIN cipher[20]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal2 ;
        RECT 83.850000 0.000000 83.920000 0.070000 ;
    END
  END cipher[20]
  PIN cipher[19]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal2 ;
        RECT 85.750000 0.000000 85.820000 0.070000 ;
    END
  END cipher[19]
  PIN cipher[18]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal2 ;
        RECT 87.650000 0.000000 87.720000 0.070000 ;
    END
  END cipher[18]
  PIN cipher[17]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal2 ;
        RECT 89.550000 0.000000 89.620000 0.070000 ;
    END
  END cipher[17]
  PIN cipher[16]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal2 ;
        RECT 91.450000 0.000000 91.520000 0.070000 ;
    END
  END cipher[16]
  PIN cipher[15]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal2 ;
        RECT 93.350000 0.000000 93.420000 0.070000 ;
    END
  END cipher[15]
  PIN cipher[14]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal2 ;
        RECT 95.250000 0.000000 95.320000 0.070000 ;
    END
  END cipher[14]
  PIN cipher[13]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal2 ;
        RECT 97.150000 0.000000 97.220000 0.070000 ;
    END
  END cipher[13]
  PIN cipher[12]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal2 ;
        RECT 99.050000 0.000000 99.120000 0.070000 ;
    END
  END cipher[12]
  PIN cipher[11]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal2 ;
        RECT 100.950000 0.000000 101.020000 0.070000 ;
    END
  END cipher[11]
  PIN cipher[10]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal2 ;
        RECT 102.850000 0.000000 102.920000 0.070000 ;
    END
  END cipher[10]
  PIN cipher[9]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal2 ;
        RECT 104.750000 0.000000 104.820000 0.070000 ;
    END
  END cipher[9]
  PIN cipher[8]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal2 ;
        RECT 106.650000 0.000000 106.720000 0.070000 ;
    END
  END cipher[8]
  PIN cipher[7]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal2 ;
        RECT 108.550000 0.000000 108.620000 0.070000 ;
    END
  END cipher[7]
  PIN cipher[6]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal2 ;
        RECT 110.450000 0.000000 110.520000 0.070000 ;
    END
  END cipher[6]
  PIN cipher[5]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal2 ;
        RECT 112.350000 0.000000 112.420000 0.070000 ;
    END
  END cipher[5]
  PIN cipher[4]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal2 ;
        RECT 114.250000 0.000000 114.320000 0.070000 ;
    END
  END cipher[4]
  PIN cipher[3]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal2 ;
        RECT 116.150000 0.000000 116.220000 0.070000 ;
    END
  END cipher[3]
  PIN cipher[2]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal2 ;
        RECT 118.050000 0.000000 118.120000 0.070000 ;
    END
  END cipher[2]
  PIN cipher[1]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal2 ;
        RECT 119.950000 0.000000 120.020000 0.070000 ;
    END
  END cipher[1]
  PIN cipher[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal2 ;
        RECT 121.850000 0.000000 121.920000 0.070000 ;
    END
  END cipher[0]
  PIN mr
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal2 ;
        RECT 91.640000 183.050000 91.710000 183.120000 ;
    END
  END mr
  PIN mw
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal2 ;
        RECT 92.590000 183.050000 92.660000 183.120000 ;
    END
  END mw
  PIN keyOrPlain[31]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal2 ;
        RECT 122.990000 183.050000 123.060000 183.120000 ;
    END
  END keyOrPlain[31]
  PIN keyOrPlain[30]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal2 ;
        RECT 122.040000 183.050000 122.110000 183.120000 ;
    END
  END keyOrPlain[30]
  PIN keyOrPlain[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal2 ;
        RECT 121.090000 183.050000 121.160000 183.120000 ;
    END
  END keyOrPlain[29]
  PIN keyOrPlain[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal2 ;
        RECT 120.140000 183.050000 120.210000 183.120000 ;
    END
  END keyOrPlain[28]
  PIN keyOrPlain[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal2 ;
        RECT 119.190000 183.050000 119.260000 183.120000 ;
    END
  END keyOrPlain[27]
  PIN keyOrPlain[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal2 ;
        RECT 118.240000 183.050000 118.310000 183.120000 ;
    END
  END keyOrPlain[26]
  PIN keyOrPlain[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal2 ;
        RECT 117.290000 183.050000 117.360000 183.120000 ;
    END
  END keyOrPlain[25]
  PIN keyOrPlain[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal2 ;
        RECT 116.340000 183.050000 116.410000 183.120000 ;
    END
  END keyOrPlain[24]
  PIN keyOrPlain[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal2 ;
        RECT 115.390000 183.050000 115.460000 183.120000 ;
    END
  END keyOrPlain[23]
  PIN keyOrPlain[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal2 ;
        RECT 114.440000 183.050000 114.510000 183.120000 ;
    END
  END keyOrPlain[22]
  PIN keyOrPlain[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal2 ;
        RECT 113.490000 183.050000 113.560000 183.120000 ;
    END
  END keyOrPlain[21]
  PIN keyOrPlain[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal2 ;
        RECT 112.540000 183.050000 112.610000 183.120000 ;
    END
  END keyOrPlain[20]
  PIN keyOrPlain[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal2 ;
        RECT 111.590000 183.050000 111.660000 183.120000 ;
    END
  END keyOrPlain[19]
  PIN keyOrPlain[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal2 ;
        RECT 110.640000 183.050000 110.710000 183.120000 ;
    END
  END keyOrPlain[18]
  PIN keyOrPlain[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal2 ;
        RECT 109.690000 183.050000 109.760000 183.120000 ;
    END
  END keyOrPlain[17]
  PIN keyOrPlain[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal2 ;
        RECT 108.740000 183.050000 108.810000 183.120000 ;
    END
  END keyOrPlain[16]
  PIN keyOrPlain[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal2 ;
        RECT 107.790000 183.050000 107.860000 183.120000 ;
    END
  END keyOrPlain[15]
  PIN keyOrPlain[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal2 ;
        RECT 106.840000 183.050000 106.910000 183.120000 ;
    END
  END keyOrPlain[14]
  PIN keyOrPlain[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal2 ;
        RECT 105.890000 183.050000 105.960000 183.120000 ;
    END
  END keyOrPlain[13]
  PIN keyOrPlain[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal2 ;
        RECT 104.940000 183.050000 105.010000 183.120000 ;
    END
  END keyOrPlain[12]
  PIN keyOrPlain[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal2 ;
        RECT 103.990000 183.050000 104.060000 183.120000 ;
    END
  END keyOrPlain[11]
  PIN keyOrPlain[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal2 ;
        RECT 103.040000 183.050000 103.110000 183.120000 ;
    END
  END keyOrPlain[10]
  PIN keyOrPlain[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal2 ;
        RECT 102.090000 183.050000 102.160000 183.120000 ;
    END
  END keyOrPlain[9]
  PIN keyOrPlain[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal2 ;
        RECT 101.140000 183.050000 101.210000 183.120000 ;
    END
  END keyOrPlain[8]
  PIN keyOrPlain[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal2 ;
        RECT 100.190000 183.050000 100.260000 183.120000 ;
    END
  END keyOrPlain[7]
  PIN keyOrPlain[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal2 ;
        RECT 99.240000 183.050000 99.310000 183.120000 ;
    END
  END keyOrPlain[6]
  PIN keyOrPlain[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal2 ;
        RECT 98.290000 183.050000 98.360000 183.120000 ;
    END
  END keyOrPlain[5]
  PIN keyOrPlain[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal2 ;
        RECT 97.340000 183.050000 97.410000 183.120000 ;
    END
  END keyOrPlain[4]
  PIN keyOrPlain[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal2 ;
        RECT 96.390000 183.050000 96.460000 183.120000 ;
    END
  END keyOrPlain[3]
  PIN keyOrPlain[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal2 ;
        RECT 95.440000 183.050000 95.510000 183.120000 ;
    END
  END keyOrPlain[2]
  PIN keyOrPlain[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal2 ;
        RECT 94.490000 183.050000 94.560000 183.120000 ;
    END
  END keyOrPlain[1]
  PIN keyOrPlain[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal2 ;
        RECT 93.540000 183.050000 93.610000 183.120000 ;
    END
  END keyOrPlain[0]
  OBS
    LAYER metal1 ;
      RECT 0.000000 0.000000 184.680000 183.120000 ;
    LAYER metal2 ;
      RECT 123.130000 182.980000 184.680000 183.120000 ;
      RECT 122.180000 182.980000 122.920000 183.120000 ;
      RECT 121.230000 182.980000 121.970000 183.120000 ;
      RECT 120.280000 182.980000 121.020000 183.120000 ;
      RECT 119.330000 182.980000 120.070000 183.120000 ;
      RECT 118.380000 182.980000 119.120000 183.120000 ;
      RECT 117.430000 182.980000 118.170000 183.120000 ;
      RECT 116.480000 182.980000 117.220000 183.120000 ;
      RECT 115.530000 182.980000 116.270000 183.120000 ;
      RECT 114.580000 182.980000 115.320000 183.120000 ;
      RECT 113.630000 182.980000 114.370000 183.120000 ;
      RECT 112.680000 182.980000 113.420000 183.120000 ;
      RECT 111.730000 182.980000 112.470000 183.120000 ;
      RECT 110.780000 182.980000 111.520000 183.120000 ;
      RECT 109.830000 182.980000 110.570000 183.120000 ;
      RECT 108.880000 182.980000 109.620000 183.120000 ;
      RECT 107.930000 182.980000 108.670000 183.120000 ;
      RECT 106.980000 182.980000 107.720000 183.120000 ;
      RECT 106.030000 182.980000 106.770000 183.120000 ;
      RECT 105.080000 182.980000 105.820000 183.120000 ;
      RECT 104.130000 182.980000 104.870000 183.120000 ;
      RECT 103.180000 182.980000 103.920000 183.120000 ;
      RECT 102.230000 182.980000 102.970000 183.120000 ;
      RECT 101.280000 182.980000 102.020000 183.120000 ;
      RECT 100.330000 182.980000 101.070000 183.120000 ;
      RECT 99.380000 182.980000 100.120000 183.120000 ;
      RECT 98.430000 182.980000 99.170000 183.120000 ;
      RECT 97.480000 182.980000 98.220000 183.120000 ;
      RECT 96.530000 182.980000 97.270000 183.120000 ;
      RECT 95.580000 182.980000 96.320000 183.120000 ;
      RECT 94.630000 182.980000 95.370000 183.120000 ;
      RECT 93.680000 182.980000 94.420000 183.120000 ;
      RECT 92.730000 182.980000 93.470000 183.120000 ;
      RECT 91.780000 182.980000 92.520000 183.120000 ;
      RECT 90.830000 182.980000 91.570000 183.120000 ;
      RECT 89.880000 182.980000 90.620000 183.120000 ;
      RECT 88.930000 182.980000 89.670000 183.120000 ;
      RECT 87.980000 182.980000 88.720000 183.120000 ;
      RECT 87.030000 182.980000 87.770000 183.120000 ;
      RECT 86.080000 182.980000 86.820000 183.120000 ;
      RECT 85.130000 182.980000 85.870000 183.120000 ;
      RECT 84.180000 182.980000 84.920000 183.120000 ;
      RECT 83.230000 182.980000 83.970000 183.120000 ;
      RECT 82.280000 182.980000 83.020000 183.120000 ;
      RECT 81.330000 182.980000 82.070000 183.120000 ;
      RECT 80.380000 182.980000 81.120000 183.120000 ;
      RECT 79.430000 182.980000 80.170000 183.120000 ;
      RECT 78.480000 182.980000 79.220000 183.120000 ;
      RECT 77.530000 182.980000 78.270000 183.120000 ;
      RECT 76.580000 182.980000 77.320000 183.120000 ;
      RECT 75.630000 182.980000 76.370000 183.120000 ;
      RECT 74.680000 182.980000 75.420000 183.120000 ;
      RECT 73.730000 182.980000 74.470000 183.120000 ;
      RECT 72.780000 182.980000 73.520000 183.120000 ;
      RECT 71.830000 182.980000 72.570000 183.120000 ;
      RECT 70.880000 182.980000 71.620000 183.120000 ;
      RECT 69.930000 182.980000 70.670000 183.120000 ;
      RECT 68.980000 182.980000 69.720000 183.120000 ;
      RECT 68.030000 182.980000 68.770000 183.120000 ;
      RECT 67.080000 182.980000 67.820000 183.120000 ;
      RECT 66.130000 182.980000 66.870000 183.120000 ;
      RECT 65.180000 182.980000 65.920000 183.120000 ;
      RECT 64.230000 182.980000 64.970000 183.120000 ;
      RECT 63.280000 182.980000 64.020000 183.120000 ;
      RECT 62.330000 182.980000 63.070000 183.120000 ;
      RECT 61.380000 182.980000 62.120000 183.120000 ;
      RECT 0.000000 182.980000 61.170000 183.120000 ;
      RECT 0.000000 0.140000 184.680000 182.980000 ;
      RECT 121.990000 0.000000 184.680000 0.140000 ;
      RECT 120.090000 0.000000 121.780000 0.140000 ;
      RECT 118.190000 0.000000 119.880000 0.140000 ;
      RECT 116.290000 0.000000 117.980000 0.140000 ;
      RECT 114.390000 0.000000 116.080000 0.140000 ;
      RECT 112.490000 0.000000 114.180000 0.140000 ;
      RECT 110.590000 0.000000 112.280000 0.140000 ;
      RECT 108.690000 0.000000 110.380000 0.140000 ;
      RECT 106.790000 0.000000 108.480000 0.140000 ;
      RECT 104.890000 0.000000 106.580000 0.140000 ;
      RECT 102.990000 0.000000 104.680000 0.140000 ;
      RECT 101.090000 0.000000 102.780000 0.140000 ;
      RECT 99.190000 0.000000 100.880000 0.140000 ;
      RECT 97.290000 0.000000 98.980000 0.140000 ;
      RECT 95.390000 0.000000 97.080000 0.140000 ;
      RECT 93.490000 0.000000 95.180000 0.140000 ;
      RECT 91.590000 0.000000 93.280000 0.140000 ;
      RECT 89.690000 0.000000 91.380000 0.140000 ;
      RECT 87.790000 0.000000 89.480000 0.140000 ;
      RECT 85.890000 0.000000 87.580000 0.140000 ;
      RECT 83.990000 0.000000 85.680000 0.140000 ;
      RECT 82.090000 0.000000 83.780000 0.140000 ;
      RECT 80.190000 0.000000 81.880000 0.140000 ;
      RECT 78.290000 0.000000 79.980000 0.140000 ;
      RECT 76.390000 0.000000 78.080000 0.140000 ;
      RECT 74.490000 0.000000 76.180000 0.140000 ;
      RECT 72.590000 0.000000 74.280000 0.140000 ;
      RECT 70.690000 0.000000 72.380000 0.140000 ;
      RECT 68.790000 0.000000 70.480000 0.140000 ;
      RECT 66.890000 0.000000 68.580000 0.140000 ;
      RECT 64.990000 0.000000 66.680000 0.140000 ;
      RECT 63.090000 0.000000 64.780000 0.140000 ;
      RECT 0.000000 0.000000 62.880000 0.140000 ;
    LAYER metal3 ;
      RECT 0.000000 0.000000 184.680000 183.120000 ;
    LAYER metal4 ;
      RECT 0.000000 0.000000 184.680000 183.120000 ;
    LAYER metal5 ;
      RECT 0.000000 0.000000 184.680000 183.120000 ;
    LAYER metal6 ;
      RECT 0.000000 0.000000 184.680000 183.120000 ;
    LAYER metal7 ;
      RECT 0.000000 0.000000 184.680000 183.120000 ;
    LAYER metal8 ;
      RECT 0.000000 0.000000 184.680000 183.120000 ;
    LAYER metal9 ;
      RECT 0.000000 0.000000 184.680000 183.120000 ;
    LAYER metal10 ;
      RECT 0.000000 0.000000 184.680000 183.120000 ;
  END
END aes128keyWrapper

END LIBRARY
