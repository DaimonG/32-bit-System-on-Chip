/ensc/cmc_homedirs/escmc29/ensc450/ENSC450finalproject/Part1/vhdl/SRAM_Lib/SRAM.lef