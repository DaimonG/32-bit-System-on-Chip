/ensc/cmc_homedirs/escmc29/ensc450/ENSC450finalproject/Part2/BE_045/results/aes128keyWrapper.lef